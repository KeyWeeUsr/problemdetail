module problemdetail

type ContentType = string

pub const type_json = 'application/problem+json'
pub const type_xml = 'application/problem+xml'
